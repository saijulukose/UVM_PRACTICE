`include "uvm_macros.svh"
import uvm_pkg::*;


module tb;
initial begin
`uvm_info("A1", "First RTL:Counter", UVM_NONE);
end

endmodule